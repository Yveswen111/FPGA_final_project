//
//
//
//

`define NM1 32'd220 //A-_freq 6-
`define NM2 32'd247 //B-_freq 7-
`define NM3 32'd262 //C_freq 1
`define NM4 32'd294 //D_freq 2
`define NM5 32'd330 //E_freq 3
`define NM6 32'd349 //F_freq 4
`define NM7 32'd392 //G_freq 5
`define NM8 32'd440 //A_freq 6
`define NM9 32'd494 //B_freq 7
`define NM10 32'd208 //G_freq+ +5-
`define NM11 32'd196 //G-_freq 5-
`define NM12 32'd524 //C+_freq 1+
`define NM13 32'd698 //F_freq+
`define NM14 32'd784 //G_freq+
`define NM15 32'd880 //A_freq+
`define NM16 32'd988 //B_freq+
`define NM15 32'd1048 //C_freq++

`define NM0 32'd20000 //slience (over freq.)

module Music (
	input [9:0] ibeatNum,	
	output reg [31:0] tone
);

always @(*) begin
	case (ibeatNum)		// 1/4 beat
		8'd0 : tone = `NM1;	//6-
		8'd1 : tone = `NM1;
		8'd2 : tone = `NM2; //7-
		8'd3 : tone = `NM2;
		8'd4 : tone = `NM3;	//1
		8'd5 : tone = `NM3;
		8'd6 : tone = `NM4; //2
		8'd7 : tone = `NM4;
		8'd8 : tone = `NM5;	//3
		8'd9 : tone = `NM5;
		8'd10 : tone = `NM5;
		8'd11 : tone = `NM5;
		8'd12 : tone = `NM8; //6
		8'd13 : tone = `NM8;
		8'd14 : tone = `NM7; //5
		8'd15 : tone = `NM7;
		8'd16 : tone = `NM5; //3
		8'd17 : tone = `NM5;
		8'd18 : tone = `NM5;
		8'd19 : tone = `NM5;
		8'd20 : tone = `NM1; //6-
		8'd21 : tone = `NM1;
		8'd22 : tone = `NM1;
		8'd23 : tone = `NM1;
		8'd24 : tone = `NM5; //3
		8'd25 : tone = `NM5;
		8'd26 : tone = `NM4; //2
		8'd27 : tone = `NM4;
		8'd28 : tone = `NM3; //1
		8'd29 : tone = `NM3;
		8'd30 : tone = `NM2; //7-
		8'd31 : tone = `NM2;
		8'd32 : tone = `NM1; //6-
		8'd33 : tone = `NM1;
		8'd34 : tone = `NM2; //7-
		8'd35 : tone = `NM2;
		8'd36 : tone = `NM3; //1
		8'd37 : tone = `NM3;
		8'd38 : tone = `NM4; //2
		8'd39 : tone = `NM4;
		8'd40 : tone = `NM5; //3
		8'd41 : tone = `NM5;
		8'd42 : tone = `NM5;
		8'd43 : tone = `NM5;
		8'd44 : tone = `NM4; //2
		8'd45 : tone = `NM4;
		8'd46 : tone = `NM3; //1
		8'd47 : tone = `NM3;
		8'd48 : tone = `NM2; //7-
		8'd49 : tone = `NM2;
		8'd50 : tone = `NM1; //6-
		8'd51 : tone = `NM1;
		8'd52 : tone = `NM2; //7-
		8'd53 : tone = `NM2;
		8'd54 : tone = `NM3; //1
		8'd55 : tone = `NM3;
		8'd56 : tone = `NM2; //7-
		8'd57 : tone = `NM2;
		8'd58 : tone = `NM1; //6-
		8'd59 : tone = `NM1;
		8'd60 : tone = `NM10; //+5-
		8'd61 : tone = `NM10;
		8'd62 : tone = `NM2; //7-
		8'd63 : tone = `NM2;
		8'd64 : tone = `NM1;//repeat
		8'd65 : tone = `NM1;
		8'd66 : tone = `NM2;
		8'd67 : tone = `NM2;
		8'd68 : tone = `NM3;
		8'd69 : tone = `NM3;
		8'd70 : tone = `NM4;
		8'd71 : tone = `NM4;
		8'd72 : tone = `NM5;
		8'd73 : tone = `NM5;
		8'd74 : tone = `NM5;
		8'd75 : tone = `NM5;
		8'd76 : tone = `NM8;
		8'd77 : tone = `NM8;
		8'd78 : tone = `NM7;
		8'd79 : tone = `NM7;
		8'd80 : tone = `NM5;
		8'd81 : tone = `NM5;
		8'd82 : tone = `NM5;
		8'd83 : tone = `NM5;
		8'd84 : tone = `NM1;
		8'd85 : tone = `NM1;
		8'd86 : tone = `NM1;
		8'd87 : tone = `NM1;
		8'd88 : tone = `NM5;
		8'd89 : tone = `NM5;
		8'd90 : tone = `NM4;
		8'd91 : tone = `NM4;
		8'd92 : tone = `NM3;
		8'd93 : tone = `NM3;
		8'd94 : tone = `NM2;
		8'd95 : tone = `NM2;
		8'd96 : tone = `NM1;
		8'd97 : tone = `NM1;
		8'd98 : tone = `NM2;
		8'd99 : tone = `NM2;
		8'd100 : tone = `NM3;
		8'd101 : tone = `NM3;
		8'd102 : tone = `NM4;
		8'd103 : tone = `NM4;
		8'd104 : tone = `NM5;
		8'd105 : tone = `NM5;
		8'd106 : tone = `NM5;
		8'd107 : tone = `NM5;
		8'd108 : tone = `NM4;
		8'd109 : tone = `NM4;
		8'd110 : tone = `NM3;
		8'd111 : tone = `NM3;
		8'd112 : tone = `NM2;
		8'd113 : tone = `NM2;
		8'd114 : tone = `NM2;
		8'd115 : tone = `NM2;
		8'd116 : tone = `NM3;
		8'd117 : tone = `NM3;
		8'd118 : tone = `NM3;
		8'd119 : tone = `NM3;
		8'd120 : tone = `NM4;
		8'd121 : tone = `NM4;
		8'd122 : tone = `NM4;
		8'd123 : tone = `NM4;
		8'd124 : tone = `NM5;
		8'd125 : tone = `NM5;
		8'd126 : tone = `NM5;
		8'd127 : tone = `NM5;
		
		
		8'd128 : tone = `NM1;	//6-
		8'd129 : tone = `NM1;
		8'd130 : tone = `NM2; //7-
		8'd131 : tone = `NM2;
		8'd132 : tone = `NM3;	//1
		8'd133 : tone = `NM3;
		8'd134 : tone = `NM4; //2
		8'd135 : tone = `NM4;
		8'd136 : tone = `NM5;	//3
		8'd137 : tone = `NM5;
		8'd138 : tone = `NM5;
		8'd139 : tone = `NM5;
		8'd140 : tone = `NM8; //6
		8'd141 : tone = `NM8;
		8'd142 : tone = `NM7; //5
		8'd143 : tone = `NM7;
		8'd144 : tone = `NM5; //3
		8'd145 : tone = `NM5;
		8'd146 : tone = `NM5;
		8'd147 : tone = `NM5;
		8'd148 : tone = `NM1; //6-
		8'd149 : tone = `NM1;
		8'd150 : tone = `NM1;
		8'd151 : tone = `NM1;
		8'd152 : tone = `NM5; //3
		8'd153 : tone = `NM5;
		8'd154 : tone = `NM4; //2
		8'd155 : tone = `NM4;
		8'd156 : tone = `NM3; //1
		8'd157 : tone = `NM3;
		8'd158 : tone = `NM2; //7-
		8'd159 : tone = `NM2;
		8'd160 : tone = `NM1; //6-
		8'd161 : tone = `NM1;
		8'd162 : tone = `NM2; //7-
		8'd163 : tone = `NM2;
		8'd164 : tone = `NM3; //1
		8'd165 : tone = `NM3;
		8'd166 : tone = `NM4; //2
		8'd167 : tone = `NM4;
		8'd168 : tone = `NM5; //3
		8'd169 : tone = `NM5;
		8'd170 : tone = `NM5;
		8'd171 : tone = `NM5;
		8'd172 : tone = `NM4; //2
		8'd173 : tone = `NM4;
		8'd174 : tone = `NM3; //1
		8'd175 : tone = `NM3;
		8'd176 : tone = `NM2; //7-
		8'd177 : tone = `NM2;
		8'd178 : tone = `NM1; //6-
		8'd179 : tone = `NM1;
		8'd180 : tone = `NM2; //7-
		8'd181 : tone = `NM2;
		8'd182 : tone = `NM3; //1
		8'd183 : tone = `NM3;
		8'd184 : tone = `NM2; //7-
		8'd185 : tone = `NM2;
		8'd186 : tone = `NM1; //6-
		8'd187 : tone = `NM1;
		8'd188 : tone = `NM10; //+5-
		8'd189 : tone = `NM10;
		8'd190 : tone = `NM2; //7-
		8'd191 : tone = `NM2;
		8'd192 : tone = `NM1;//repeat
		8'd193 : tone = `NM1;
		8'd194 : tone = `NM2;
		8'd195 : tone = `NM2;
		8'd196 : tone = `NM3;
		8'd197 : tone = `NM3;
		8'd198 : tone = `NM4;
		8'd199 : tone = `NM4;
		8'd200 : tone = `NM5;
		8'd201 : tone = `NM5;
		8'd202 : tone = `NM5;
		8'd203 : tone = `NM5;
		8'd204 : tone = `NM8;
		8'd205 : tone = `NM8;
		8'd206 : tone = `NM7;
		8'd207 : tone = `NM7;
		8'd208 : tone = `NM5;
		8'd209 : tone = `NM5;
		8'd210 : tone = `NM5;
		8'd211 : tone = `NM5;
		8'd212 : tone = `NM1;
		8'd213 : tone = `NM1;
		8'd214 : tone = `NM1;
		8'd215 : tone = `NM1;
		8'd216 : tone = `NM5;
		8'd217 : tone = `NM5;
		8'd218 : tone = `NM4;
		8'd219 : tone = `NM4;
		8'd220 : tone = `NM3;
		8'd221 : tone = `NM3;
		8'd222 : tone = `NM2;
		8'd223 : tone = `NM2;
		8'd224 : tone = `NM1;
		8'd225 : tone = `NM1;
		8'd226 : tone = `NM2;
		8'd227 : tone = `NM2;
		8'd228 : tone = `NM3;
		8'd229 : tone = `NM3;
		8'd230 : tone = `NM4;
		8'd231 : tone = `NM4;
		8'd232 : tone = `NM5;
		8'd233 : tone = `NM5;
		8'd234 : tone = `NM5;
		8'd235 : tone = `NM5;
		8'd236 : tone = `NM4;
		8'd237 : tone = `NM4;
		8'd238 : tone = `NM3;
		8'd239 : tone = `NM3;
		8'd240 : tone = `NM2;
		8'd241 : tone = `NM2;
		8'd242 : tone = `NM2;
		8'd243 : tone = `NM2;
		8'd244 : tone = `NM3;
		8'd245 : tone = `NM3;
		8'd246 : tone = `NM3;
		8'd247 : tone = `NM3;
		8'd248 : tone = `NM4;
		8'd249 : tone = `NM4;
		8'd250 : tone = `NM4;
		8'd251 : tone = `NM4;
		8'd252 : tone = `NM5;
		8'd253 : tone = `NM5;
		8'd254 : tone = `NM5;
		8'd255 : tone = `NM5;
		
		8'd256 : tone = `NM7;
		8'd257 : tone = `NM7;
		8'd258 : tone = `NM8;
		8'd259 : tone = `NM8;
		8'd260 : tone = `NM5;
		8'd261 : tone = `NM5;
		8'd262 : tone = `NM4;
		8'd263 : tone = `NM4;
		8'd264 : tone = `NM5;
		8'd265 : tone = `NM5;
		8'd266 : tone = `NM5;
		8'd267 : tone = `NM5;
		8'd268 : tone = `NM4;
		8'd269 : tone = `NM4;
		8'd270 : tone = `NM5;
		8'd271 : tone = `NM5;
		
		8'd272 : tone = `NM7;
		8'd273 : tone = `NM7;
		8'd274 : tone = `NM8;
		8'd275 : tone = `NM8;
		8'd276 : tone = `NM5;
		8'd277 : tone = `NM5;
		8'd278 : tone = `NM4;
		8'd279 : tone = `NM4;
		8'd280 : tone = `NM5;
		8'd281 : tone = `NM5;
		8'd282 : tone = `NM5;
		8'd283 : tone = `NM5;
		8'd284 : tone = `NM4;
		8'd285 : tone = `NM4;
		8'd286 : tone = `NM5;
		8'd287 : tone = `NM5;
		
		8'd288 : tone = `NM4;
		8'd289 : tone = `NM4;
		8'd290 : tone = `NM3;
		8'd291 : tone = `NM3;
		8'd292 : tone = `NM2;
		8'd293 : tone = `NM2;
		8'd294 : tone = `NM11;
		8'd295 : tone = `NM11;
		8'd296 : tone = `NM1;
		8'd297 : tone = `NM1;
		8'd298 : tone = `NM1;
		8'd299 : tone = `NM1;
		8'd300 : tone = `NM11;
		8'd301 : tone = `NM11;
		8'd302 : tone = `NM1;
		8'd303 : tone = `NM1;
		
		8'd304 : tone = `NM2;
		8'd305 : tone = `NM2;
		8'd306 : tone = `NM3;
		8'd307 : tone = `NM3;
		8'd308 : tone = `NM4;
		8'd309 : tone = `NM4;
		8'd310 : tone = `NM5;
		8'd311 : tone = `NM5;
		8'd312 : tone = `NM1;
		8'd313 : tone = `NM1;
		8'd314 : tone = `NM1;
		8'd315 : tone = `NM1;
		8'd316 : tone = `NM5;
		8'd317 : tone = `NM5;
		8'd318 : tone = `NM7;
		8'd319 : tone = `NM7;
		
		8'd320 : tone = `NM7;
		8'd321 : tone = `NM7;
		8'd322 : tone = `NM8;
		8'd323 : tone = `NM8;
		8'd324 : tone = `NM5;
		8'd325 : tone = `NM5;
		8'd326 : tone = `NM4;
		8'd327 : tone = `NM4;
		8'd328 : tone = `NM5;
		8'd329 : tone = `NM5;
		8'd330 : tone = `NM5;
		8'd331 : tone = `NM5;
		8'd332 : tone = `NM4;
		8'd333 : tone = `NM4;
		8'd334 : tone = `NM5;
		8'd335 : tone = `NM5;
		
		8'd336 : tone = `NM7;
		8'd337 : tone = `NM7;
		8'd338 : tone = `NM8;
		8'd339 : tone = `NM8;
		8'd340 : tone = `NM5;
		8'd341 : tone = `NM5;
		8'd342 : tone = `NM4;
		8'd343 : tone = `NM4;
		8'd344 : tone = `NM5;
		8'd345 : tone = `NM5;
		8'd346 : tone = `NM5;
		8'd347 : tone = `NM5;
		8'd348 : tone = `NM4;
		8'd349 : tone = `NM4;
		8'd350 : tone = `NM5;
		8'd351 : tone = `NM5;
		
		8'd352 : tone = `NM4;
		8'd353 : tone = `NM4;
		8'd354 : tone = `NM3;
		8'd355 : tone = `NM3;
		8'd356 : tone = `NM2;
		8'd357 : tone = `NM2;
		8'd358 : tone = `NM11;
		8'd359 : tone = `NM11;
		8'd360 : tone = `NM1;
		8'd361 : tone = `NM1;
		8'd362 : tone = `NM1;
		8'd363 : tone = `NM1;
		8'd364 : tone = `NM11;
		8'd365 : tone = `NM11;
		8'd366 : tone = `NM1;
		8'd367 : tone = `NM1;
		
		8'd368 : tone = `NM2;
		8'd369 : tone = `NM2;
		8'd370 : tone = `NM3;
		8'd371 : tone = `NM3;
		8'd372 : tone = `NM4;
		8'd373 : tone = `NM4;
		8'd374 : tone = `NM5;
		8'd375 : tone = `NM5;
		8'd376 : tone = `NM1;
		8'd377 : tone = `NM1;
		8'd378 : tone = `NM1;
		8'd379 : tone = `NM1;
		8'd380 : tone = `NM5;
		8'd381 : tone = `NM5;
		8'd382 : tone = `NM7;
		8'd383 : tone = `NM7;
	
		8'd384 : tone = `NM7;
		8'd385 : tone = `NM7;
		8'd386 : tone = `NM8;
		8'd387 : tone = `NM8;
		8'd388 : tone = `NM5;
		8'd389 : tone = `NM5;
		8'd390 : tone = `NM4;
		8'd391 : tone = `NM4;
		8'd392 : tone = `NM5;
		8'd393 : tone = `NM5;
		8'd394 : tone = `NM5;
		8'd395 : tone = `NM5;
		8'd396 : tone = `NM4;
		8'd397 : tone = `NM4;
		8'd398 : tone = `NM5;
		8'd399 : tone = `NM5;
		
		8'd400 : tone = `NM7;
		8'd401 : tone = `NM7;
		8'd402 : tone = `NM8;
		8'd403 : tone = `NM8;
		8'd404 : tone = `NM5;
		8'd405 : tone = `NM5;
		8'd406 : tone = `NM4;
		8'd407 : tone = `NM4;
		8'd408 : tone = `NM5;
		8'd409 : tone = `NM5;
		8'd410 : tone = `NM5;
		8'd411 : tone = `NM5;
		8'd412 : tone = `NM4;
		8'd413 : tone = `NM4;
		8'd414 : tone = `NM5;
		8'd415 : tone = `NM5;

		8'd416 : tone = `NM4;
		8'd417 : tone = `NM4;
		8'd418 : tone = `NM3;
		8'd419 : tone = `NM3;
		8'd420 : tone = `NM2;
		8'd421 : tone = `NM2;
		8'd422 : tone = `NM11;
		8'd423 : tone = `NM11;
		8'd424 : tone = `NM1;
		8'd425 : tone = `NM1;
		8'd426 : tone = `NM1;
		8'd427 : tone = `NM1;
		8'd428 : tone = `NM11;
		8'd429 : tone = `NM11;
		8'd430 : tone = `NM1;
		8'd431 : tone = `NM1;

		8'd432 : tone = `NM2;
		8'd433 : tone = `NM2;
		8'd434 : tone = `NM3;
		8'd435 : tone = `NM3;
		8'd436 : tone = `NM4;
		8'd437 : tone = `NM4;
		8'd438 : tone = `NM5;
		8'd439 : tone = `NM5;
		8'd440 : tone = `NM1;
		8'd441 : tone = `NM1;
		8'd442 : tone = `NM1;
		8'd443 : tone = `NM1;
		8'd444 : tone = `NM5;
		8'd445 : tone = `NM5;
		8'd446 : tone = `NM7;
		8'd447 : tone = `NM7;
		
		8'd448 : tone = `NM7;
		8'd449 : tone = `NM7;
		8'd450 : tone = `NM8;
		8'd451 : tone = `NM8;
		8'd452 : tone = `NM5;
		8'd453 : tone = `NM5;
		8'd454 : tone = `NM4;
		8'd455 : tone = `NM4;
		8'd456 : tone = `NM5;
		8'd457 : tone = `NM5;
		8'd458 : tone = `NM5;
		8'd459 : tone = `NM5;
		8'd460 : tone = `NM4;
		8'd461 : tone = `NM4;
		8'd462 : tone = `NM5;
		8'd463 : tone = `NM5;
		
		8'd464 : tone = `NM7;
		8'd465 : tone = `NM7;
		8'd466 : tone = `NM8;
		8'd467 : tone = `NM8;
		8'd468 : tone = `NM5;
		8'd469 : tone = `NM5;
		8'd470 : tone = `NM4;
		8'd471 : tone = `NM4;
		8'd472 : tone = `NM5;
		8'd473 : tone = `NM5;
		8'd474 : tone = `NM5;
		8'd475 : tone = `NM5;
		8'd476 : tone = `NM8;
		8'd477 : tone = `NM8;
		8'd478 : tone = `NM9;
		8'd479 : tone = `NM9;

		8'd480 : tone = `NM12;
		8'd481 : tone = `NM12;
		8'd482 : tone = `NM9;
		8'd483 : tone = `NM9;
		8'd484 : tone = `NM8;
		8'd485 : tone = `NM8;
		8'd486 : tone = `NM7;
		8'd487 : tone = `NM7;
		8'd488 : tone = `NM5;
		8'd489 : tone = `NM5;
		8'd490 : tone = `NM5;
		8'd491 : tone = `NM5;
		8'd492 : tone = `NM4;
		8'd493 : tone = `NM4;
		8'd494 : tone = `NM5;
		8'd495 : tone = `NM5;

		8'd496 : tone = `NM4;
		8'd497 : tone = `NM4;
		8'd498 : tone = `NM3;
		8'd499 : tone = `NM3;
		8'd500 : tone = `NM2;
		8'd501 : tone = `NM2;
		8'd502 : tone = `NM11;
		8'd503 : tone = `NM11;
		8'd504 : tone = `NM1;
		8'd505 : tone = `NM1;
		8'd506 : tone = `NM1;
		8'd507 : tone = `NM1;
		8'd508 : tone = `NM5;
		8'd509 : tone = `NM5;
		8'd510 : tone = `NM7;
		8'd511 : tone = `NM7;
		
		8'd512 : tone = `NM7;
		8'd513 : tone = `NM7;
		8'd514 : tone = `NM8;
		8'd515 : tone = `NM8;
		8'd516 : tone = `NM5;
		8'd517 : tone = `NM5;
		8'd518 : tone = `NM4;
		8'd519 : tone = `NM4;
		8'd520 : tone = `NM5;
		8'd521 : tone = `NM5;
		8'd522 : tone = `NM5;
		8'd523 : tone = `NM5;
		8'd524 : tone = `NM4;
		8'd525 : tone = `NM4;
		8'd526 : tone = `NM5;
		8'd527 : tone = `NM5;
		
		8'd528 : tone = `NM7;
		8'd529 : tone = `NM7;
		8'd530 : tone = `NM8;
		8'd531 : tone = `NM8;
		8'd532 : tone = `NM5;
		8'd533 : tone = `NM5;
		8'd534 : tone = `NM4;
		8'd535 : tone = `NM4;
		8'd536 : tone = `NM5;
		8'd537 : tone = `NM5;
		8'd538 : tone = `NM5;
		8'd539 : tone = `NM5;
		8'd540 : tone = `NM4;
		8'd541 : tone = `NM4;
		8'd542 : tone = `NM5;
		8'd543 : tone = `NM5;

		8'd544 : tone = `NM4;
		8'd545 : tone = `NM4;
		8'd546 : tone = `NM3;
		8'd547 : tone = `NM3;
		8'd548 : tone = `NM2;
		8'd549 : tone = `NM2;
		8'd550 : tone = `NM11;
		8'd551 : tone = `NM11;
		8'd552 : tone = `NM1;
		8'd553 : tone = `NM1;
		8'd554 : tone = `NM1;
		8'd555 : tone = `NM1;
		8'd556 : tone = `NM11;
		8'd557 : tone = `NM11;
		8'd558 : tone = `NM1;
		8'd559 : tone = `NM1;

		8'd560 : tone = `NM2;
		8'd561 : tone = `NM2;
		8'd562 : tone = `NM3;
		8'd563 : tone = `NM3;
		8'd564 : tone = `NM4;
		8'd565 : tone = `NM4;
		8'd567 : tone = `NM5;
		8'd568 : tone = `NM5;
		8'd569 : tone = `NM1;
		8'd570 : tone = `NM1;
		8'd571 : tone = `NM1;
		8'd572 : tone = `NM1;
		8'd573 : tone = `NM5;
		8'd574 : tone = `NM5;
		8'd575 : tone = `NM7;
		8'd576 : tone = `NM7;
	
		8'd577 : tone = `NM7;
		8'd578 : tone = `NM7;
		8'd579 : tone = `NM8;
		8'd580 : tone = `NM8;
		8'd581 : tone = `NM5;
		8'd582 : tone = `NM5;
		8'd583 : tone = `NM4;
		8'd584 : tone = `NM4;
		8'd585 : tone = `NM5;
		8'd586 : tone = `NM5;
		8'd587 : tone = `NM5;
		8'd588 : tone = `NM5;
		8'd589 : tone = `NM4;
		8'd590 : tone = `NM4;
		8'd591 : tone = `NM5;
		8'd592 : tone = `NM5;

		8'd593 : tone = `NM7;
		8'd594 : tone = `NM7;
		8'd595 : tone = `NM8;
		8'd596 : tone = `NM8;
		8'd597 : tone = `NM5;
		8'd598 : tone = `NM5;
		8'd599 : tone = `NM4;
		8'd600 : tone = `NM4;
		8'd601 : tone = `NM5;
		8'd602 : tone = `NM5;
		8'd603 : tone = `NM5;
		8'd604 : tone = `NM5;
		8'd605 : tone = `NM4;
		8'd606 : tone = `NM4;
		8'd607 : tone = `NM5;
		8'd608 : tone = `NM5;
	
		8'd609 : tone = `NM4;
		8'd610 : tone = `NM4;
		8'd611 : tone = `NM3;
		8'd612 : tone = `NM3;
		8'd613 : tone = `NM2;
		8'd614 : tone = `NM2;
		8'd615 : tone = `NM11;
		8'd616 : tone = `NM11;
		8'd617 : tone = `NM1;
		8'd618 : tone = `NM1;
		8'd619 : tone = `NM1;
		8'd620 : tone = `NM1;
		8'd621 : tone = `NM11;
		8'd622 : tone = `NM11;
		8'd623 : tone = `NM1;
		8'd624 : tone = `NM1;

		8'd625 : tone = `NM2;
		8'd626 : tone = `NM2;
		8'd627 : tone = `NM3;
		8'd628 : tone = `NM3;
		8'd629 : tone = `NM4;
		8'd630 : tone = `NM4;
		8'd631 : tone = `NM5;
		8'd632 : tone = `NM5;
		8'd633 : tone = `NM1;
		8'd634 : tone = `NM1;
		8'd635 : tone = `NM1;
		8'd636 : tone = `NM1;
		8'd637 : tone = `NM5;
		8'd638 : tone = `NM5;
		8'd639 : tone = `NM7;
		8'd640 : tone = `NM7;

		8'd641 : tone = `NM7;
		8'd642 : tone = `NM7;
		8'd643 : tone = `NM8;
		8'd644 : tone = `NM8;
		8'd645 : tone = `NM5;
		8'd646 : tone = `NM5;
		8'd647 : tone = `NM4;
		8'd648 : tone = `NM4;
		8'd649 : tone = `NM5;
		8'd650 : tone = `NM5;
		8'd651 : tone = `NM5;
		8'd652 : tone = `NM5;
		8'd653 : tone = `NM4;
		8'd654 : tone = `NM4;
		8'd655 : tone = `NM5;
		8'd656 : tone = `NM5;
	
		8'd657 : tone = `NM7;
		8'd658 : tone = `NM7;
		8'd659 : tone = `NM8;
		8'd660 : tone = `NM8;
		8'd661 : tone = `NM5;
		8'd662 : tone = `NM5;
		8'd663 : tone = `NM4;
		8'd664 : tone = `NM4;
		8'd665 : tone = `NM5;
		8'd666 : tone = `NM5;
		8'd667 : tone = `NM5;
		8'd668 : tone = `NM5;
		8'd669 : tone = `NM4;
		8'd670 : tone = `NM4;
		8'd671 : tone = `NM5;
		8'd672 : tone = `NM5;
		
		8'd673 : tone = `NM4;
		8'd674 : tone = `NM4;
		8'd675 : tone = `NM3;
		8'd676 : tone = `NM3;
		8'd677 : tone = `NM2;
		8'd678 : tone = `NM2;
		8'd679 : tone = `NM11;
		8'd680 : tone = `NM11;
		8'd681 : tone = `NM1;
		8'd682 : tone = `NM1;
		8'd683 : tone = `NM1;
		8'd684 : tone = `NM1;
		8'd685 : tone = `NM11;
		8'd686 : tone = `NM11;
		8'd687 : tone = `NM1;
		8'd688 : tone = `NM1;
		
		8'd689 : tone = `NM2;
		8'd690 : tone = `NM2;
		8'd691 : tone = `NM3;
		8'd692 : tone = `NM3;
		8'd693 : tone = `NM4;
		8'd694 : tone = `NM4;
		8'd695 : tone = `NM5;
		8'd696 : tone = `NM5;
		8'd697 : tone = `NM1;
		8'd698 : tone = `NM1;
		8'd699 : tone = `NM1;
		8'd700 : tone = `NM1;
		8'd701 : tone = `NM5;
		8'd702 : tone = `NM5;
		8'd703 : tone = `NM7;
		8'd704 : tone = `NM7;
	
		8'd705 : tone = `NM7;
		8'd706 : tone = `NM7;
		8'd707 : tone = `NM8;
		8'd708 : tone = `NM8;
		8'd709 : tone = `NM5;
		8'd710 : tone = `NM5;
		8'd711 : tone = `NM4;
		8'd712 : tone = `NM4;
		8'd713 : tone = `NM5;
		8'd714 : tone = `NM5;
		8'd715 : tone = `NM5;
		8'd716 : tone = `NM5;
		8'd717 : tone = `NM4;
		8'd718 : tone = `NM4;
		8'd719 : tone = `NM5;
		8'd720 : tone = `NM5;
	
		8'd721 : tone = `NM7;
		8'd722 : tone = `NM7;
		8'd723 : tone = `NM8;
		8'd724 : tone = `NM8;
		8'd725 : tone = `NM5;
		8'd726 : tone = `NM5;
		8'd727 : tone = `NM4;
		8'd728 : tone = `NM4;
		8'd729 : tone = `NM5;
		8'd730 : tone = `NM5;
		8'd731 : tone = `NM5;
		8'd732 : tone = `NM5;
		8'd733 : tone = `NM8;
		8'd734 : tone = `NM8;
		8'd735 : tone = `NM9;
		8'd736 : tone = `NM9;
		
		8'd737 : tone = `NM12;
		8'd738 : tone = `NM12;
		8'd739 : tone = `NM9;
		8'd740 : tone = `NM9;
		8'd741 : tone = `NM8;
		8'd742 : tone = `NM8;
		8'd743 : tone = `NM7;
		8'd744 : tone = `NM7;
		8'd745 : tone = `NM5;
		8'd746 : tone = `NM5;
		8'd747 : tone = `NM5;
		8'd748 : tone = `NM5;
		8'd749 : tone = `NM4;
		8'd750 : tone = `NM4;
		8'd751 : tone = `NM5;
		8'd752 : tone = `NM5;
		
		8'd753 : tone = `NM4;
		8'd754 : tone = `NM4;
		8'd755 : tone = `NM3;
		8'd756 : tone = `NM3;
		8'd757 : tone = `NM2;
		8'd758 : tone = `NM2;
		8'd759 : tone = `NM11;
		8'd760 : tone = `NM11;
		8'd761 : tone = `NM1;
		8'd762 : tone = `NM1;
		8'd763 : tone = `NM1;
		8'd764 : tone = `NM1;
		8'd765 : tone = `NM0;
		8'd766 : tone = `NM0;
		8'd767 : tone = `NM0;
		8'd768 : tone = `NM0;
		
		default : tone = `NM0;
	endcase
end

endmodule