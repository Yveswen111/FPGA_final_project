`define NM1 32'd220 //A-_freq 6-
`define NM2 32'd247 //B-_freq 7-
`define NM3 32'd262 //C_freq 1
`define NM4 32'd294 //D_freq 2
`define NM5 32'd330 //E_freq 3
`define NM6 32'd349 //F_freq 4
`define NM7 32'd392 //G_freq 5
`define NM8 32'd440 //A_freq 6
`define NM9 32'd494 //B_freq 7
`define NM10 32'd208 //G_freq+ +5-
`define NM11 32'd196 //G-_freq 5-
`define NM12 32'd524 //C+_freq 1+
`define NM13 32'd698 //F_freq+
`define NM14 32'd784 //G_freq+
`define NM15 32'd880 //A_freq+
`define NM16 32'd988 //B_freq+
`define NM17 32'd1048 //C_freq++

`define NM0 32'd20000 //slience (over freq.)

module Music_game (
	input [9:0] ibeatNum,	
	output reg [31:0] tone
);

always @(*) begin
	case (ibeatNum)		// 1/4 beat
		10'd0 : tone = `NM1;	//6-
		10'd1 : tone = `NM1;
		10'd2 : tone = `NM2; //7-
		10'd3 : tone = `NM2;
		10'd4 : tone = `NM3;	//1
		10'd5 : tone = `NM3;
		10'd6 : tone = `NM4; //2
		10'd7 : tone = `NM4;
		10'd8 : tone = `NM5;	//3
		10'd9 : tone = `NM5;
		10'd10 : tone = `NM5;
		10'd11 : tone = `NM5;
		10'd12 : tone = `NM8; //6
		10'd13 : tone = `NM8;
		10'd14 : tone = `NM7; //5
		10'd15 : tone = `NM7;
		10'd16 : tone = `NM5; //3
		10'd17 : tone = `NM5;
		10'd18 : tone = `NM5;
		10'd19 : tone = `NM5;
		10'd20 : tone = `NM1; //6-
		10'd21 : tone = `NM1;
		10'd22 : tone = `NM1;
		10'd23 : tone = `NM1;
		10'd24 : tone = `NM5; //3
		10'd25 : tone = `NM5;
		10'd26 : tone = `NM4; //2
		10'd27 : tone = `NM4;
		10'd28 : tone = `NM3; //1
		10'd29 : tone = `NM3;
		10'd30 : tone = `NM2; //7-
		10'd31 : tone = `NM2;
		10'd32 : tone = `NM1; //6-
		10'd33 : tone = `NM1;
		10'd34 : tone = `NM2; //7-
		10'd35 : tone = `NM2;
		10'd36 : tone = `NM3; //1
		10'd37 : tone = `NM3;
		10'd38 : tone = `NM4; //2
		10'd39 : tone = `NM4;
		10'd40 : tone = `NM5; //3
		10'd41 : tone = `NM5;
		10'd42 : tone = `NM5;
		10'd43 : tone = `NM5;
		10'd44 : tone = `NM4; //2
		10'd45 : tone = `NM4;
		10'd46 : tone = `NM3; //1
		10'd47 : tone = `NM3;
		10'd48 : tone = `NM2; //7-
		10'd49 : tone = `NM2;
		10'd50 : tone = `NM1; //6-
		10'd51 : tone = `NM1;
		10'd52 : tone = `NM2; //7-
		10'd53 : tone = `NM2;
		10'd54 : tone = `NM3; //1
		10'd55 : tone = `NM3;
		10'd56 : tone = `NM2; //7-
		10'd57 : tone = `NM2;
		10'd58 : tone = `NM1; //6-
		10'd59 : tone = `NM1;
		10'd60 : tone = `NM10; //+5-
		10'd61 : tone = `NM10;
		10'd62 : tone = `NM2; //7-
		10'd63 : tone = `NM2;
		10'd64 : tone = `NM1;//repeat
		10'd65 : tone = `NM1;
		10'd66 : tone = `NM2;
		10'd67 : tone = `NM2;
		10'd68 : tone = `NM3;
		10'd69 : tone = `NM3;
		10'd70 : tone = `NM4;
		10'd71 : tone = `NM4;
		10'd72 : tone = `NM5;
		10'd73 : tone = `NM5;
		10'd74 : tone = `NM5;
		10'd75 : tone = `NM5;
		10'd76 : tone = `NM8;
		10'd77 : tone = `NM8;
		10'd78 : tone = `NM7;
		10'd79 : tone = `NM7;
		10'd80 : tone = `NM5;
		10'd81 : tone = `NM5;
		10'd82 : tone = `NM5;
		10'd83 : tone = `NM5;
		10'd84 : tone = `NM1;
		10'd85 : tone = `NM1;
		10'd86 : tone = `NM1;
		10'd87 : tone = `NM1;
		10'd88 : tone = `NM5;
		10'd89 : tone = `NM5;
		10'd90 : tone = `NM4;
		10'd91 : tone = `NM4;
		10'd92 : tone = `NM3;
		10'd93 : tone = `NM3;
		10'd94 : tone = `NM2;
		10'd95 : tone = `NM2;
		10'd96 : tone = `NM1;
		10'd97 : tone = `NM1;
		10'd98 : tone = `NM2;
		10'd99 : tone = `NM2;
		10'd100 : tone = `NM3;
		10'd101 : tone = `NM3;
		10'd102 : tone = `NM4;
		10'd103 : tone = `NM4;
		10'd104 : tone = `NM5;
		10'd105 : tone = `NM5;
		10'd106 : tone = `NM5;
		10'd107 : tone = `NM5;
		10'd108 : tone = `NM4;
		10'd109 : tone = `NM4;
		10'd110 : tone = `NM3;
		10'd111 : tone = `NM3;
		10'd112 : tone = `NM2;
		10'd113 : tone = `NM2;
		10'd114 : tone = `NM2;
		10'd115 : tone = `NM2;
		10'd116 : tone = `NM3;
		10'd117 : tone = `NM3;
		10'd118 : tone = `NM3;
		10'd119 : tone = `NM3;
		10'd120 : tone = `NM4;
		10'd121 : tone = `NM4;
		10'd122 : tone = `NM4;
		10'd123 : tone = `NM4;
		10'd124 : tone = `NM5;
		10'd125 : tone = `NM5;
		10'd126 : tone = `NM5;
		10'd127 : tone = `NM5;
		
		
		10'd128 : tone = `NM1;	//6-
		10'd129 : tone = `NM1;
		10'd130 : tone = `NM2; //7-
		10'd131 : tone = `NM2;
		10'd132 : tone = `NM3;	//1
		10'd133 : tone = `NM3;
		10'd134 : tone = `NM4; //2
		10'd135 : tone = `NM4;
		10'd136 : tone = `NM5;	//3
		10'd137 : tone = `NM5;
		10'd138 : tone = `NM5;
		10'd139 : tone = `NM5;
		10'd140 : tone = `NM8; //6
		10'd141 : tone = `NM8;
		10'd142 : tone = `NM7; //5
		10'd143 : tone = `NM7;
		10'd144 : tone = `NM5; //3
		10'd145 : tone = `NM5;
		10'd146 : tone = `NM5;
		10'd147 : tone = `NM5;
		10'd148 : tone = `NM1; //6-
		10'd149 : tone = `NM1;
		10'd150 : tone = `NM1;
		10'd151 : tone = `NM1;
		10'd152 : tone = `NM5; //3
		10'd153 : tone = `NM5;
		10'd154 : tone = `NM4; //2
		10'd155 : tone = `NM4;
		10'd156 : tone = `NM3; //1
		10'd157 : tone = `NM3;
		10'd158 : tone = `NM2; //7-
		10'd159 : tone = `NM2;
		10'd160 : tone = `NM1; //6-
		10'd161 : tone = `NM1;
		10'd162 : tone = `NM2; //7-
		10'd163 : tone = `NM2;
		10'd164 : tone = `NM3; //1
		10'd165 : tone = `NM3;
		10'd166 : tone = `NM4; //2
		10'd167 : tone = `NM4;
		10'd168 : tone = `NM5; //3
		10'd169 : tone = `NM5;
		10'd170 : tone = `NM5;
		10'd171 : tone = `NM5;
		10'd172 : tone = `NM4; //2
		10'd173 : tone = `NM4;
		10'd174 : tone = `NM3; //1
		10'd175 : tone = `NM3;
		10'd176 : tone = `NM2; //7-
		10'd177 : tone = `NM2;
		10'd178 : tone = `NM1; //6-
		10'd179 : tone = `NM1;
		10'd180 : tone = `NM2; //7-
		10'd181 : tone = `NM2;
		10'd182 : tone = `NM3; //1
		10'd183 : tone = `NM3;
		10'd184 : tone = `NM2; //7-
		10'd185 : tone = `NM2;
		10'd186 : tone = `NM1; //6-
		10'd187 : tone = `NM1;
		10'd188 : tone = `NM10; //+5-
		10'd189 : tone = `NM10;
		10'd190 : tone = `NM2; //7-
		10'd191 : tone = `NM2;
		10'd192 : tone = `NM1;//repeat
		10'd193 : tone = `NM1;
		10'd194 : tone = `NM2;
		10'd195 : tone = `NM2;
		10'd196 : tone = `NM3;
		10'd197 : tone = `NM3;
		10'd198 : tone = `NM4;
		10'd199 : tone = `NM4;
		10'd200 : tone = `NM5;
		10'd201 : tone = `NM5;
		10'd202 : tone = `NM5;
		10'd203 : tone = `NM5;
		10'd204 : tone = `NM8;
		10'd205 : tone = `NM8;
		10'd206 : tone = `NM7;
		10'd207 : tone = `NM7;
		10'd208 : tone = `NM5;
		10'd209 : tone = `NM5;
		10'd210 : tone = `NM5;
		10'd211 : tone = `NM5;
		10'd212 : tone = `NM1;
		10'd213 : tone = `NM1;
		10'd214 : tone = `NM1;
		10'd215 : tone = `NM1;
		10'd216 : tone = `NM5;
		10'd217 : tone = `NM5;
		10'd218 : tone = `NM4;
		10'd219 : tone = `NM4;
		10'd220 : tone = `NM3;
		10'd221 : tone = `NM3;
		10'd222 : tone = `NM2;
		10'd223 : tone = `NM2;
		10'd224 : tone = `NM1;
		10'd225 : tone = `NM1;
		10'd226 : tone = `NM2;
		10'd227 : tone = `NM2;
		10'd228 : tone = `NM3;
		10'd229 : tone = `NM3;
		10'd230 : tone = `NM4;
		10'd231 : tone = `NM4;
		10'd232 : tone = `NM5;
		10'd233 : tone = `NM5;
		10'd234 : tone = `NM5;
		10'd235 : tone = `NM5;
		10'd236 : tone = `NM4;
		10'd237 : tone = `NM4;
		10'd238 : tone = `NM3;
		10'd239 : tone = `NM3;
		10'd240 : tone = `NM2;
		10'd241 : tone = `NM2;
		10'd242 : tone = `NM2;
		10'd243 : tone = `NM2;
		10'd244 : tone = `NM3;
		10'd245 : tone = `NM3;
		10'd246 : tone = `NM3;
		10'd247 : tone = `NM3;
		10'd248 : tone = `NM4;
		10'd249 : tone = `NM4;
		10'd250 : tone = `NM4;
		10'd251 : tone = `NM4;
		10'd252 : tone = `NM5;
		10'd253 : tone = `NM5;
		10'd254 : tone = `NM5;
		10'd255 : tone = `NM5;
		
		10'd256 : tone = `NM7;
		10'd257 : tone = `NM7;
		10'd258 : tone = `NM8;
		10'd259 : tone = `NM8;
		10'd260 : tone = `NM5;
		10'd261 : tone = `NM5;
		10'd262 : tone = `NM4;
		10'd263 : tone = `NM4;
		10'd264 : tone = `NM5;
		10'd265 : tone = `NM5;
		10'd266 : tone = `NM5;
		10'd267 : tone = `NM5;
		10'd268 : tone = `NM4;
		10'd269 : tone = `NM4;
		10'd270 : tone = `NM5;
		10'd271 : tone = `NM5;
		
		10'd272 : tone = `NM7;
		10'd273 : tone = `NM7;
		10'd274 : tone = `NM8;
		10'd275 : tone = `NM8;
		10'd276 : tone = `NM5;
		10'd277 : tone = `NM5;
		10'd278 : tone = `NM4;
		10'd279 : tone = `NM4;
		10'd280 : tone = `NM5;
		10'd281 : tone = `NM5;
		10'd282 : tone = `NM5;
		10'd283 : tone = `NM5;
		10'd284 : tone = `NM4;
		10'd285 : tone = `NM4;
		10'd286 : tone = `NM5;
		10'd287 : tone = `NM5;
		
		10'd288 : tone = `NM4;
		10'd289 : tone = `NM4;
		10'd290 : tone = `NM3;
		10'd291 : tone = `NM3;
		10'd292 : tone = `NM2;
		10'd293 : tone = `NM2;
		10'd294 : tone = `NM11;
		10'd295 : tone = `NM11;
		10'd296 : tone = `NM1;
		10'd297 : tone = `NM1;
		10'd298 : tone = `NM1;
		10'd299 : tone = `NM1;
		10'd300 : tone = `NM11;
		10'd301 : tone = `NM11;
		10'd302 : tone = `NM1;
		10'd303 : tone = `NM1;
		
		10'd304 : tone = `NM2;
		10'd305 : tone = `NM2;
		10'd306 : tone = `NM3;
		10'd307 : tone = `NM3;
		10'd308 : tone = `NM4;
		10'd309 : tone = `NM4;
		10'd310 : tone = `NM5;
		10'd311 : tone = `NM5;
		10'd312 : tone = `NM1;
		10'd313 : tone = `NM1;
		10'd314 : tone = `NM1;
		10'd315 : tone = `NM1;
		10'd316 : tone = `NM5;
		10'd317 : tone = `NM5;
		10'd318 : tone = `NM7;
		10'd319 : tone = `NM7;
		
		10'd320 : tone = `NM7;
		10'd321 : tone = `NM7;
		10'd322 : tone = `NM8;
		10'd323 : tone = `NM8;
		10'd324 : tone = `NM5;
		10'd325 : tone = `NM5;
		10'd326 : tone = `NM4;
		10'd327 : tone = `NM4;
		10'd328 : tone = `NM5;
		10'd329 : tone = `NM5;
		10'd330 : tone = `NM5;
		10'd331 : tone = `NM5;
		10'd332 : tone = `NM4;
		10'd333 : tone = `NM4;
		10'd334 : tone = `NM5;
		10'd335 : tone = `NM5;
		
		10'd336 : tone = `NM7;
		10'd337 : tone = `NM7;
		10'd338 : tone = `NM8;
		10'd339 : tone = `NM8;
		10'd340 : tone = `NM5;
		10'd341 : tone = `NM5;
		10'd342 : tone = `NM4;
		10'd343 : tone = `NM4;
		10'd344 : tone = `NM5;
		10'd345 : tone = `NM5;
		10'd346 : tone = `NM5;
		10'd347 : tone = `NM5;
		10'd348 : tone = `NM4;
		10'd349 : tone = `NM4;
		10'd350 : tone = `NM5;
		10'd351 : tone = `NM5;
		
		10'd352 : tone = `NM4;
		10'd353 : tone = `NM4;
		10'd354 : tone = `NM3;
		10'd355 : tone = `NM3;
		10'd356 : tone = `NM2;
		10'd357 : tone = `NM2;
		10'd358 : tone = `NM11;
		10'd359 : tone = `NM11;
		10'd360 : tone = `NM1;
		10'd361 : tone = `NM1;
		10'd362 : tone = `NM1;
		10'd363 : tone = `NM1;
		10'd364 : tone = `NM11;
		10'd365 : tone = `NM11;
		10'd366 : tone = `NM1;
		10'd367 : tone = `NM1;
		
		10'd368 : tone = `NM2;
		10'd369 : tone = `NM2;
		10'd370 : tone = `NM3;
		10'd371 : tone = `NM3;
		10'd372 : tone = `NM4;
		10'd373 : tone = `NM4;
		10'd374 : tone = `NM5;
		10'd375 : tone = `NM5;
		10'd376 : tone = `NM1;
		10'd377 : tone = `NM1;
		10'd378 : tone = `NM1;
		10'd379 : tone = `NM1;
		10'd380 : tone = `NM5;
		10'd381 : tone = `NM5;
		10'd382 : tone = `NM7;
		10'd383 : tone = `NM7;
	
		10'd384 : tone = `NM7;
		10'd385 : tone = `NM7;
		10'd386 : tone = `NM8;
		10'd387 : tone = `NM8;
		10'd388 : tone = `NM5;
		10'd389 : tone = `NM5;
		10'd390 : tone = `NM4;
		10'd391 : tone = `NM4;
		10'd392 : tone = `NM5;
		10'd393 : tone = `NM5;
		10'd394 : tone = `NM5;
		10'd395 : tone = `NM5;
		10'd396 : tone = `NM4;
		10'd397 : tone = `NM4;
		10'd398 : tone = `NM5;
		10'd399 : tone = `NM5;
		
		10'd400 : tone = `NM7;
		10'd401 : tone = `NM7;
		10'd402 : tone = `NM8;
		10'd403 : tone = `NM8;
		10'd404 : tone = `NM5;
		10'd405 : tone = `NM5;
		10'd406 : tone = `NM4;
		10'd407 : tone = `NM4;
		10'd408 : tone = `NM5;
		10'd409 : tone = `NM5;
		10'd410 : tone = `NM5;
		10'd411 : tone = `NM5;
		10'd412 : tone = `NM4;
		10'd413 : tone = `NM4;
		10'd414 : tone = `NM5;
		10'd415 : tone = `NM5;

		10'd416 : tone = `NM4;
		10'd417 : tone = `NM4;
		10'd418 : tone = `NM3;
		10'd419 : tone = `NM3;
		10'd420 : tone = `NM2;
		10'd421 : tone = `NM2;
		10'd422 : tone = `NM11;
		10'd423 : tone = `NM11;
		10'd424 : tone = `NM1;
		10'd425 : tone = `NM1;
		10'd426 : tone = `NM1;
		10'd427 : tone = `NM1;
		10'd428 : tone = `NM11;
		10'd429 : tone = `NM11;
		10'd430 : tone = `NM1;
		10'd431 : tone = `NM1;

		10'd432 : tone = `NM2;
		10'd433 : tone = `NM2;
		10'd434 : tone = `NM3;
		10'd435 : tone = `NM3;
		10'd436 : tone = `NM4;
		10'd437 : tone = `NM4;
		10'd438 : tone = `NM5;
		10'd439 : tone = `NM5;
		10'd440 : tone = `NM1;
		10'd441 : tone = `NM1;
		10'd442 : tone = `NM1;
		10'd443 : tone = `NM1;
		10'd444 : tone = `NM5;
		10'd445 : tone = `NM5;
		10'd446 : tone = `NM7;
		10'd447 : tone = `NM7;
		
		10'd448 : tone = `NM7;
		10'd449 : tone = `NM7;
		10'd450 : tone = `NM8;
		10'd451 : tone = `NM8;
		10'd452 : tone = `NM5;
		10'd453 : tone = `NM5;
		10'd454 : tone = `NM4;
		10'd455 : tone = `NM4;
		10'd456 : tone = `NM5;
		10'd457 : tone = `NM5;
		10'd458 : tone = `NM5;
		10'd459 : tone = `NM5;
		10'd460 : tone = `NM4;
		10'd461 : tone = `NM4;
		10'd462 : tone = `NM5;
		10'd463 : tone = `NM5;
		
		10'd464 : tone = `NM7;
		10'd465 : tone = `NM7;
		10'd466 : tone = `NM8;
		10'd467 : tone = `NM8;
		10'd468 : tone = `NM5;
		10'd469 : tone = `NM5;
		10'd470 : tone = `NM4;
		10'd471 : tone = `NM4;
		10'd472 : tone = `NM5;
		10'd473 : tone = `NM5;
		10'd474 : tone = `NM5;
		10'd475 : tone = `NM5;
		10'd476 : tone = `NM8;
		10'd477 : tone = `NM8;
		10'd478 : tone = `NM9;
		10'd479 : tone = `NM9;

		10'd480 : tone = `NM12;
		10'd481 : tone = `NM12;
		10'd482 : tone = `NM9;
		10'd483 : tone = `NM9;
		10'd484 : tone = `NM8;
		10'd485 : tone = `NM8;
		10'd486 : tone = `NM7;
		10'd487 : tone = `NM7;
		10'd488 : tone = `NM5;
		10'd489 : tone = `NM5;
		10'd490 : tone = `NM5;
		10'd491 : tone = `NM5;
		10'd492 : tone = `NM4;
		10'd493 : tone = `NM4;
		10'd494 : tone = `NM5;
		10'd495 : tone = `NM5;

		10'd496 : tone = `NM4;
		10'd497 : tone = `NM4;
		10'd498 : tone = `NM3;
		10'd499 : tone = `NM3;
		10'd500 : tone = `NM2;
		10'd501 : tone = `NM2;
		10'd502 : tone = `NM11;
		10'd503 : tone = `NM11;
		10'd504 : tone = `NM1;
		10'd505 : tone = `NM1;
		10'd506 : tone = `NM1;
		10'd507 : tone = `NM1;
		10'd508 : tone = `NM5;
		10'd509 : tone = `NM5;
		10'd510 : tone = `NM7;
		10'd511 : tone = `NM7;
		
		10'd512 : tone = `NM7;
		10'd513 : tone = `NM7;
		10'd514 : tone = `NM8;
		10'd515 : tone = `NM8;
		10'd516 : tone = `NM5;
		10'd517 : tone = `NM5;
		10'd518 : tone = `NM4;
		10'd519 : tone = `NM4;
		10'd520 : tone = `NM5;
		10'd521 : tone = `NM5;
		10'd522 : tone = `NM5;
		10'd523 : tone = `NM5;
		10'd524 : tone = `NM4;
		10'd525 : tone = `NM4;
		10'd526 : tone = `NM5;
		10'd527 : tone = `NM5;
		
		10'd528 : tone = `NM7;
		10'd529 : tone = `NM7;
		10'd530 : tone = `NM8;
		10'd531 : tone = `NM8;
		10'd532 : tone = `NM5;
		10'd533 : tone = `NM5;
		10'd534 : tone = `NM4;
		10'd535 : tone = `NM4;
		10'd536 : tone = `NM5;
		10'd537 : tone = `NM5;
		10'd538 : tone = `NM5;
		10'd539 : tone = `NM5;
		10'd540 : tone = `NM4;
		10'd541 : tone = `NM4;
		10'd542 : tone = `NM5;
		10'd543 : tone = `NM5;

		10'd544 : tone = `NM4;
		10'd545 : tone = `NM4;
		10'd546 : tone = `NM3;
		10'd547 : tone = `NM3;
		10'd548 : tone = `NM2;
		10'd549 : tone = `NM2;
		10'd550 : tone = `NM11;
		10'd551 : tone = `NM11;
		10'd552 : tone = `NM1;
		10'd553 : tone = `NM1;
		10'd554 : tone = `NM1;
		10'd555 : tone = `NM1;
		10'd556 : tone = `NM11;
		10'd557 : tone = `NM11;
		10'd558 : tone = `NM1;
		10'd559 : tone = `NM1;

		10'd560 : tone = `NM2;
		10'd561 : tone = `NM2;
		10'd562 : tone = `NM3;
		10'd563 : tone = `NM3;
		10'd564 : tone = `NM4;
		10'd565 : tone = `NM4;
		10'd567 : tone = `NM5;
		10'd568 : tone = `NM5;
		10'd569 : tone = `NM1;
		10'd570 : tone = `NM1;
		10'd571 : tone = `NM1;
		10'd572 : tone = `NM1;
		10'd573 : tone = `NM5;
		10'd574 : tone = `NM5;
		10'd575 : tone = `NM7;
		10'd576 : tone = `NM7;
	
		10'd577 : tone = `NM7;
		10'd578 : tone = `NM7;
		10'd579 : tone = `NM8;
		10'd580 : tone = `NM8;
		10'd581 : tone = `NM5;
		10'd582 : tone = `NM5;
		10'd583 : tone = `NM4;
		10'd584 : tone = `NM4;
		10'd585 : tone = `NM5;
		10'd586 : tone = `NM5;
		10'd587 : tone = `NM5;
		10'd588 : tone = `NM5;
		10'd589 : tone = `NM4;
		10'd590 : tone = `NM4;
		10'd591 : tone = `NM5;
		10'd592 : tone = `NM5;

		10'd593 : tone = `NM7;
		10'd594 : tone = `NM7;
		10'd595 : tone = `NM8;
		10'd596 : tone = `NM8;
		10'd597 : tone = `NM5;
		10'd598 : tone = `NM5;
		10'd599 : tone = `NM4;
		10'd600 : tone = `NM4;
		10'd601 : tone = `NM5;
		10'd602 : tone = `NM5;
		10'd603 : tone = `NM5;
		10'd604 : tone = `NM5;
		10'd605 : tone = `NM4;
		10'd606 : tone = `NM4;
		10'd607 : tone = `NM5;
		10'd608 : tone = `NM5;
	
		10'd609 : tone = `NM4;
		10'd610 : tone = `NM4;
		10'd611 : tone = `NM3;
		10'd612 : tone = `NM3;
		10'd613 : tone = `NM2;
		10'd614 : tone = `NM2;
		10'd615 : tone = `NM11;
		10'd616 : tone = `NM11;
		10'd617 : tone = `NM1;
		10'd618 : tone = `NM1;
		10'd619 : tone = `NM1;
		10'd620 : tone = `NM1;
		10'd621 : tone = `NM11;
		10'd622 : tone = `NM11;
		10'd623 : tone = `NM1;
		10'd624 : tone = `NM1;

		10'd625 : tone = `NM2;
		10'd626 : tone = `NM2;
		10'd627 : tone = `NM3;
		10'd628 : tone = `NM3;
		10'd629 : tone = `NM4;
		10'd630 : tone = `NM4;
		10'd631 : tone = `NM5;
		10'd632 : tone = `NM5;
		10'd633 : tone = `NM1;
		10'd634 : tone = `NM1;
		10'd635 : tone = `NM1;
		10'd636 : tone = `NM1;
		10'd637 : tone = `NM5;
		10'd638 : tone = `NM5;
		10'd639 : tone = `NM7;
		10'd640 : tone = `NM7;

		10'd641 : tone = `NM7;
		10'd642 : tone = `NM7;
		10'd643 : tone = `NM8;
		10'd644 : tone = `NM8;
		10'd645 : tone = `NM5;
		10'd646 : tone = `NM5;
		10'd647 : tone = `NM4;
		10'd648 : tone = `NM4;
		10'd649 : tone = `NM5;
		10'd650 : tone = `NM5;
		10'd651 : tone = `NM5;
		10'd652 : tone = `NM5;
		10'd653 : tone = `NM4;
		10'd654 : tone = `NM4;
		10'd655 : tone = `NM5;
		10'd656 : tone = `NM5;
	
		10'd657 : tone = `NM7;
		10'd658 : tone = `NM7;
		10'd659 : tone = `NM8;
		10'd660 : tone = `NM8;
		10'd661 : tone = `NM5;
		10'd662 : tone = `NM5;
		10'd663 : tone = `NM4;
		10'd664 : tone = `NM4;
		10'd665 : tone = `NM5;
		10'd666 : tone = `NM5;
		10'd667 : tone = `NM5;
		10'd668 : tone = `NM5;
		10'd669 : tone = `NM4;
		10'd670 : tone = `NM4;
		10'd671 : tone = `NM5;
		10'd672 : tone = `NM5;
		
		10'd673 : tone = `NM4;
		10'd674 : tone = `NM4;
		10'd675 : tone = `NM3;
		10'd676 : tone = `NM3;
		10'd677 : tone = `NM2;
		10'd678 : tone = `NM2;
		10'd679 : tone = `NM11;
		10'd680 : tone = `NM11;
		10'd681 : tone = `NM1;
		10'd682 : tone = `NM1;
		10'd683 : tone = `NM1;
		10'd684 : tone = `NM1;
		10'd685 : tone = `NM11;
		10'd686 : tone = `NM11;
		10'd687 : tone = `NM1;
		10'd688 : tone = `NM1;
		
		10'd689 : tone = `NM2;
		10'd690 : tone = `NM2;
		10'd691 : tone = `NM3;
		10'd692 : tone = `NM3;
		10'd693 : tone = `NM4;
		10'd694 : tone = `NM4;
		10'd695 : tone = `NM5;
		10'd696 : tone = `NM5;
		10'd697 : tone = `NM1;
		10'd698 : tone = `NM1;
		10'd699 : tone = `NM1;
		10'd700 : tone = `NM1;
		10'd701 : tone = `NM5;
		10'd702 : tone = `NM5;
		10'd703 : tone = `NM7;
		10'd704 : tone = `NM7;
	
		10'd705 : tone = `NM7;
		10'd706 : tone = `NM7;
		10'd707 : tone = `NM8;
		10'd708 : tone = `NM8;
		10'd709 : tone = `NM5;
		10'd710 : tone = `NM5;
		10'd711 : tone = `NM4;
		10'd712 : tone = `NM4;
		10'd713 : tone = `NM5;
		10'd714 : tone = `NM5;
		10'd715 : tone = `NM5;
		10'd716 : tone = `NM5;
		10'd717 : tone = `NM4;
		10'd718 : tone = `NM4;
		10'd719 : tone = `NM5;
		10'd720 : tone = `NM5;
	
		10'd721 : tone = `NM7;
		10'd722 : tone = `NM7;
		10'd723 : tone = `NM8;
		10'd724 : tone = `NM8;
		10'd725 : tone = `NM5;
		10'd726 : tone = `NM5;
		10'd727 : tone = `NM4;
		10'd728 : tone = `NM4;
		10'd729 : tone = `NM5;
		10'd730 : tone = `NM5;
		10'd731 : tone = `NM5;
		10'd732 : tone = `NM5;
		10'd733 : tone = `NM8;
		10'd734 : tone = `NM8;
		10'd735 : tone = `NM9;
		10'd736 : tone = `NM9;
		
		10'd737 : tone = `NM12;
		10'd738 : tone = `NM12;
		10'd739 : tone = `NM9;
		10'd740 : tone = `NM9;
		10'd741 : tone = `NM8;
		10'd742 : tone = `NM8;
		10'd743 : tone = `NM7;
		10'd744 : tone = `NM7;
		10'd745 : tone = `NM5;
		10'd746 : tone = `NM5;
		10'd747 : tone = `NM5;
		10'd748 : tone = `NM5;
		10'd749 : tone = `NM4;
		10'd750 : tone = `NM4;
		10'd751 : tone = `NM5;
		10'd752 : tone = `NM5;
		
		10'd753 : tone = `NM4;
		10'd754 : tone = `NM4;
		10'd755 : tone = `NM3;
		10'd756 : tone = `NM3;
		10'd757 : tone = `NM2;
		10'd758 : tone = `NM2;
		10'd759 : tone = `NM11;
		10'd760 : tone = `NM11;
		10'd761 : tone = `NM1;
		10'd762 : tone = `NM1;
		10'd763 : tone = `NM1;
		10'd764 : tone = `NM1;
		10'd765 : tone = `NM0;
		10'd766 : tone = `NM0;
		10'd767 : tone = `NM0;
		10'd768 : tone = `NM0;
		
		default : tone = `NM0;
	endcase
end

endmodule